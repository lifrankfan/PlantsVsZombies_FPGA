module pvz_background_rom (
	input logic clock,
	input logic [17:0] address,
	output logic [3:0] q
);

logic [3:0] memory [0:153599] /* synthesis ram_init_file = "./pvz_background/pvz_background.COE" */;

always_ff @ (posedge clock) begin
	q <= memory[address];
end

endmodule
